interface and_if();

logic A, B;
logic Y;

modport DUT(input A, B, output Y);
endinterface