module and_DUT(and_if.DUT intf);


assign intf.Y=intf.A & intf.B;

endmodule